netcdf ecmwf{ // European Centre for Medium-Range Weather Forecasts (ECMWF) model


dimensions:
        record = UNLIMITED ;  // (reference time, forecast time)
        lat = 73 ;            // latitude
        lon = 145 ;           // longitude
        level = 4 ;           // isobaric levels
        time_len = 21 ;       // string length for datetime strings
        valtime_offset = 9 ;  // number of offset times
        nmodels = 29 ;         // number of models
        ngrids = 12 ;         // number of grids
        nav = 1 ;             // for navigation
        nav_len = 100 ;       // max string length for navigation strings

variables:

        double reftime(record) ;	// reference time of the model
               reftime:long_name = "reference time" ;
               reftime:units = "hours since 1992-1-1" ;

        double valtime(record) ;	// forecast time ("valid" time)
               valtime:long_name = "valid time" ;
               valtime:units = "hours since 1992-1-1" ;

        :record = "reftime, valtime" ;	// "dimension attribute" -- means
                                        // (reftime, valtime) uniquely
                                        // determine record

        char   datetime(record, time_len) ; // derived from reftime
               datetime:long_name = "reference date and time" ;
               // units YYYY-MM-DD hh:mm:ssZ  (ISO 8601)

        double valtime_offset(valtime_offset) ; // valtime - reftime
               valtime_offset:long_name = "hours from reference time" ;
               valtime_offset:units = "hours" ;

        char   forecasttime(record, time_len) ; // derived from valtime
               forecasttime:long_name = "forecast date and time" ;
               // units YYYY-MM-DD hh:mm:ssZ  (ISO 8601)

        float  level(level) ;
               level:long_name = "isobaric level" ;
               level:units = "hectopascals" ;


        // The following lat and lon coordinate variables are redundant,
        // since the navigation variables provide the necessary information.
        // The extra information is included here for human readability.

        float  lat(lat) ;
               lat:long_name = "latitude" ;
               lat:units = "degrees_north" ;

        float  lon(lon) ;
               lon:long_name = "longitude" ;
               lon:units = "degrees_east" ;

        long   model_id(nmodels) ;
               model_id:long_name = "generating process ID number" ;

        // navigation variables all use nav dimension

        char   nav_model(nav, nav_len) ;        // navigation parameterization
               nav_model:long_name = "navigation model name" ;

        int    grid_type_code(nav) ;
               grid_type_code:long_name = "GRIB-1 GDS data representation type" ;

        char   grid_type(nav, nav_len) ;
               grid_type:long_name = "GRIB-1 grid type" ;

        char   grid_name(nav, nav_len) ;
               grid_name:long_name = "grid name" ;

        int    grid_center(nav) ;
               grid_center:long_name = "GRIB-1 originating center ID" ;

        int    grid_number(nav, ngrids) ;
               grid_number:long_name = "GRIB-1 catalogued grid numbers" ;
               grid_number:_FillValue = -9999 ;

        char   i_dim(nav, nav_len) ;
               i_dim:long_name = "longitude dimension name" ;

        char   j_dim(nav, nav_len) ;
               j_dim:long_name = "latitude dimension name" ;

        int    Ni(nav) ;
               Ni:long_name = "number of points along a latitude circle" ;

        int    Nj(nav) ;
               Nj:long_name = "number of points along a longitude circle" ;

        float  La1(nav) ;
               La1:long_name = "latitude of first grid point" ;
               La1:units = "degrees_north" ;

        float  Lo1(nav) ;
               Lo1:long_name = "longitude of first grid point" ;
               Lo1:units = "degrees_east" ;

        float  La2(nav) ;
               La2:long_name = "latitude of last grid point" ;
               La2:units = "degrees_north" ;

        float  Lo2(nav) ;
               Lo2:long_name = "longitude of last grid point" ;
               Lo2:units = "degrees_east" ;

        float  Di(nav) ;
               Di:long_name = "longitudinal direction increment" ;
               Di:units = "degrees" ;

        float  Dj(nav) ;
               Dj:long_name = "latitudinal direction increment" ;
               Dj:units = "degrees" ;

        byte   ResCompFlag(nav) ;
               ResCompFlag:long_name = "resolution and component flags" ;

        // end of navigation variables

        float  T(record,level,lat,lon) ;
               T:long_name = "Temperature at isobaric levels" ;
               T:standard_name = "air_temperature" ;
               T:units = "degK" ;
               T:GRIB_parameter_number = 11 ;
               T:GRIB_level_flag = 100 ;
               T:_FillValue = -9999.f ;
               T:navigation = "nav" ;

        float  RH(record,level,lat,lon) ;
               RH:long_name = "Relative humidity at isobaric levels" ;
               RH:standard_name = "relative_humidity" ;
               RH:units = "percent" ;
               RH:GRIB_parameter_number = 52 ;
               RH:GRIB_level_flag = 100 ;
               RH:_FillValue = -9999.f ;
               RH:navigation = "nav" ;

        float  P_msl_sfc(record,lat,lon) ;
               P_msl_sfc:long_name = "Pressure reduced to MSL at surface of the earth" ;
               P_msl_sfc:standard_name = "air_pressure_at_sea_level" ;
               P_msl_sfc:units = "Pa" ;
               P_msl_sfc:GRIB_parameter_number = 2 ;
               P_msl_sfc:GRIB_level_flag = 1 ;
               P_msl_sfc:_FillValue = -9999.f ;
               P_msl_sfc:navigation = "nav" ;

        float  Z(record,level,lat,lon) ;
               Z:long_name = "Geopotential height at isobaric levels" ;
               Z:standard_name = "geopotential_height" ;
               Z:units = "gp m" ;
               Z:GRIB_parameter_number = 7 ;
               Z:GRIB_level_flag = 100 ;
               Z:_FillValue = -9999.f ;
               Z:navigation = "nav" ;

        float  u(record,level,lat,lon) ;
               u:long_name = "u-component of wind at isobaric levels" ;
               u:standard_name = "eastward_wind" ;
               u:units = "m/s" ;
               u:GRIB_parameter_number = 33 ;
               u:GRIB_level_flag = 100 ;
               u:_FillValue = -9999.f ;
               u:navigation = "nav" ;

        float  v(record,level,lat,lon) ;
               v:long_name = "v-component of wind at isobaric levels" ;
               v:standard_name = "northward_wind" ;
               v:units = "m/s" ;
               v:GRIB_parameter_number = 34 ;
               v:GRIB_level_flag = 100 ;
               v:_FillValue = -9999.f ;
               v:navigation = "nav" ;


// global attributes
               :history = "2003-03-28 11:58:27 - created by gribtocdl" ; 
               :title = "European Centre for Medium-Range Weather Forecasts model" ;
               :Conventions = "NUWG" ;
               :GRIB_reference = "Office Note 388 GRIB" ;
               :GRIB_URL = "http://www.nco.ncep.noaa.gov/pmb/docs/on388/" ;
               :version = 1.0 ;

data:

 level = 850.0, 700.0, 500.0, 200.0 ;
 model_id = 202, 203, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132,
   133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147;
 valtime_offset = 0, 24, 48, 72, 96, 120, 144, 168, 204 ;


 // Navigation
 nav_model = "GRIB1" ;
 grid_type_code = 0 ;
 grid_type = "Latitude/Longitude" ;
 grid_name = "Global 5.0 x 2.5 degree grid" ;
 grid_center = 98 ;
 grid_number = 1,2,3,4,5,6,7,8,9,10,11,12 ;   // stitched together
 i_dim = "lon" ;
 j_dim = "lat" ;
 Ni = 73 ;
 Nj = 145 ;
 La1 = -90.000000 ;
 Lo1 = -180.000000 ;
 La2 = 90.000000 ;
 Lo2 = 180.000000 ;
 Di = 2.500000 ;
 Dj = 2.500000 ;
 ResCompFlag = 128 ;

 lon = -180.0,-177.5,-175.0,-172.5,-170.0,-167.5,-165.0,-162.5,
       -160.0,-157.5,-155.0,-152.5,-150.0,-147.5,-145.0,-142.5,
       -140.0,-137.5,-135.0,-132.5,-130.0,-127.5,-125.0,-122.5,
       -120.0,-117.5,-115.0,-112.5,-110.0,-107.5,-105.0,-102.5,
       -100.0, -97.5, -95.0, -92.5, -90.0, -87.5, -85.0, -82.5,
        -80.0, -77.5, -75.0, -72.5, -70.0, -67.5, -65.0, -62.5,
        -60.0, -57.5, -55.0, -52.5, -50.0, -47.5, -45.0, -42.5,
        -40.0, -37.5, -35.0, -32.5, -30.0, -27.5, -25.0, -22.5,
        -20.0, -17.5, -15.0, -12.5, -10.0,  -7.5,  -5.0,  -2.5,
          0.0,   2.5,   5.0,   7.5,  10.0,  12.5,  15.0,  17.5,
         20.0,  22.5,  25.0,  27.5,  30.0,  32.5,  35.0,  37.5,
         40.0,  42.5,  45.0,  47.5,  50.0,  52.5,  55.0,  57.5,
         60.0,  62.5,  65.0,  67.5,  70.0,  72.5,  75.0,  77.5,
         80.0,  82.5,  85.0,  87.5,  90.0,  92.5,  95.0,  97.5,
        100.0, 102.5, 105.0, 107.5, 110.0, 112.5, 115.0, 117.5,
        120.0, 122.5, 125.0, 127.5, 130.0, 132.5, 135.0, 137.5,
        140.0, 142.5, 145.0, 147.5, 150.0, 152.5, 155.0, 157.5,
        160.0, 162.5, 165.0, 167.5, 170.0, 172.5, 175.0, 177.5, 180.0 ;

 lat = -90.0,-87.5,-85.0,-82.5,-80.0,-77.5,-75.0,-72.5,
       -70.0,-67.5,-65.0,-62.5,-60.0,-57.5,-55.0,-52.5,
       -50.0,-47.5,-45.0,-42.5,-40.0,-37.5,-35.0,-32.5,
       -30.0,-27.5,-25.0,-22.5,-20.0,-17.5,-15.0,-12.5,
       -10.0, -7.5, -5.0, -2.5,  0.0,  2.5,  5.0,  7.5,
        10.0, 12.5, 15.0, 17.5, 20.0, 22.5, 25.0, 27.5,
        30.0, 32.5, 35.0, 37.5, 40.0, 42.5, 45.0, 47.5,
        50.0, 52.5, 55.0, 57.5, 60.0, 62.5, 65.0, 67.5,
        70.0, 72.5, 75.0, 77.5, 80.0, 82.5, 85.0, 87.5, 90.0 ;

}
