netcdf sst-t {          // Sea Surface Temperature Analysis Model

dimensions:
        record = UNLIMITED ;   // (reference time, forecast time)
        lat = 91 ;             // latitude
        lon = 181 ;            // longitude
        time_len = 21 ;        // string length for datetime strings
        valtime_offset = 1 ;   // number of offset times
        nmodels = 1 ;          // number of models
        ngrids = 4 ;           // number of grids
        nav = 1 ;              // for navigation
        nav_len = 100 ;        // max string length for navigation strings

variables:

        double reftime(record) ;	// reference time of the model
               reftime:long_name = "reference time" ;
               reftime:units = "hours since 1992-1-1" ;

        double valtime(record) ;	// forecast time ("valid" time)
               valtime:long_name = "valid time" ;
               valtime:units = "hours since 1992-1-1" ;

        :record = "reftime, valtime" ;	// "dimension attribute" -- means
                                        // (reftime, valtime) uniquely
                                        // determine record

        char   datetime(record, time_len) ; // derived from reftime
               datetime:long_name = "reference date and time" ;
               // units YYYY-MM-DD hh:mm:ssZ  (ISO 8601)

        double valtime_offset(valtime_offset) ; // valtime - reftime
               valtime_offset:long_name = "hours from reference time" ;
               valtime_offset:units = "hours" ;

        char   forecasttime(record, time_len) ; // derived from valtime
               forecasttime:long_name = "forecast date and time" ;
               // units YYYY-MM-DD hh:mm:ssZ  (ISO 8601)


        // The following lat and lon coordinate variables are redundant,
        // since the navigation variables provide the necessary information.
        // The extra information is included here for human readability.

        float  lat(lat) ;
               lat:long_name = "latitude" ;
               lat:units = "degrees_north" ;

        float  lon(lon) ;
               lon:long_name = "longitude" ;
               lon:units = "degrees_east" ;

        long   model_id(nmodels) ;
               model_id:long_name = "generating process ID number" ;

        // navigation variables all use nav dimension

        char   nav_model(nav, nav_len) ;        // navigation parameterization
               nav_model:long_name = "navigation model name" ;

        int    grid_type_code(nav) ;
               grid_type_code:long_name = "GRIB-1 GDS data representation type" ;

        char   grid_type(nav, nav_len) ;
               grid_type:long_name = "GRIB-1 grid type" ;

        char   grid_name(nav, nav_len) ;
               grid_name:long_name = "grid name" ;

        int    grid_center(nav) ;
               grid_center:long_name = "GRIB-1 originating center ID" ;

        int    grid_number(nav, ngrids) ;
               grid_number:long_name = "GRIB-1 catalogued grid numbers" ;
               grid_number:_FillValue = -9999 ;

        char   i_dim(nav, nav_len) ;
               i_dim:long_name = "longitude dimension name" ;

        char   j_dim(nav, nav_len) ;
               j_dim:long_name = "latitude dimension name" ;

        int    Ni(nav) ;
               Ni:long_name = "number of points along a latitude circle" ;

        int    Nj(nav) ;
               Nj:long_name = "number of points along a longitude circle" ;

        float  La1(nav) ;
               La1:long_name = "latitude of first grid point" ;
               La1:units = "degrees_north" ;

        float  Lo1(nav) ;
               Lo1:long_name = "longitude of first grid point" ;
               Lo1:units = "degrees_east" ;

        float  La2(nav) ;
               La2:long_name = "latitude of last grid point" ;
               La2:units = "degrees_north" ;

        float  Lo2(nav) ;
               Lo2:long_name = "longitude of last grid point" ;
               Lo2:units = "degrees_east" ;

        float  Di(nav) ;
               Di:long_name = "longitudinal direction increment" ;
               Di:units = "degrees" ;

        float  Dj(nav) ;
               Dj:long_name = "latitudinal direction increment" ;
               Dj:units = "degrees" ;

        byte   ResCompFlag(nav) ;
               ResCompFlag:long_name = "resolution and component flags" ;

        // end of navigation variables

        float  SST(record, lat, lon) ;
               SST:long_name = "Sea temperature" ;
               SST:standard_name = "sea_water_temperature" ;
               SST:units = "degK" ;
               SST:GRIB_parameter_number = 80 ;
               SST:GRIB_level_flag = 1 ;
               SST:_FillValue = -9999.f ;
               SST:navigation = "nav" ;

// global attributes
               :history = "2003-04-07 12:12:50 - created by gribtocdl" ; 
               :title = "Sea Surface Temperature Analysis Model" ;
               :Conventions = "NUWG" ;
               :GRIB_reference = "Office Note 388 GRIB" ;
               :GRIB_URL = "http://www.nco.ncep.noaa.gov/pmb/docs/on388/" ;
               :version = 1.0 ;

data:

 model_id = 44 ;
 valtime_offset = 0 ;


 // Navigation
 nav_model = "GRIB1" ;
 grid_type_code = 0 ;
 grid_type = "Latitude/Longitude" ;
 grid_name = "Global 2.0 x 2.0 degree grid" ;
 grid_center = 7 ;  // NCEP
 grid_number = 61, 62, 63, 64 ;
 i_dim = "lon" ;
 j_dim = "lat" ;
 Ni = 181 ;
 Nj = 91 ;
 La1 = -90.000000 ;
 Lo1 = -180.000000 ;
 La2 = 90.000000 ;
 Lo2 = 180.000000 ;
 Di = 2.000000 ;
 Dj = 2.000000 ;
 ResCompFlag = 136 ;

 lon = -180,-178,-176,-174,-172,-170,-168,-166,-164,-162,
       -160,-158,-156,-154,-152,-150,-148,-146,-144,-142,
       -140,-138,-136,-134,-132,-130,-128,-126,-124,-122,
       -120,-118,-116,-114,-112,-110,-108,-106,-104,-102,
       -100, -98, -96, -94, -92, -90, -88, -86, -84, -82,
        -80, -78, -76, -74, -72, -70, -68, -66, -64, -62,
        -60, -58, -56, -54, -52, -50, -48, -46, -44, -42,
        -40, -38, -36, -34, -32, -30, -28, -26, -24, -22,
        -20, -18, -16, -14, -12, -10,  -8,  -6,  -4,  -2,
          0,   2,   4,   6,   8,  10,  12,  14,  16,  18,
         20,  22,  24,  26,  28,  30,  32,  34,  36,  38,
         40,  42,  44,  46,  48,  50,  52,  54,  56,  58,
         60,  62,  64,  66,  68,  70,  72,  74,  76,  78,
         80,  82,  84,  86,  88,  90,  92,  94,  96,  98,
        100, 102, 104, 106, 108, 110, 112, 114, 116, 118,
        120, 122, 124, 126, 128, 130, 132, 134, 136, 138,
        140, 142, 144, 146, 148, 150, 152, 154, 156, 158,
        160, 162, 164, 166, 168, 170, 172, 174, 176, 178, 180 ;

 lat = -90,-88,-86,-84,-82,-80,-78,-76,-74,-72,-70,-68,-66,-64,-62,
       -60,-58,-56,-54,-52,-50,-48,-46,-44,-42,-40,-38,-36,-34,-32,
       -30,-28,-26,-24,-22,-20,-18,-16,-14,-12,-10, -8, -6, -4, -2,
         0,  2,  4,  6,  8, 10, 12, 14, 16, 18, 20, 22, 24, 26, 28,
        30, 32, 34, 36, 38, 40, 42, 44, 46, 48, 50, 52, 54, 56, 58,
        60, 62, 64, 66, 68, 70, 72, 74, 76, 78, 80, 82, 84, 86, 88, 90 ;

}
