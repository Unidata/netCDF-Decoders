netcdf mrf-e{            // Medium Range Forecasts Extended


dimensions:
        record = UNLIMITED ;  // (reference time, forecast time)
        lat = 37 ;            // latitude
        lon = 72 ;            // longitude
        level = 2 ;           // isobaric levels
        time_len = 21 ;       // string length for datetime strings
        valtime_offset = 14 ; // number of offset times
        nmodels = 2 ;         // number of models
        ngrids = 2 ;          // number of grids
        nav = 1 ;             // for navigation
        nav_len = 100 ;       // max string length for navigation strings

variables:

        double reftime(record) ;	// reference time of the model
               reftime:long_name = "reference time" ;
               reftime:units = "hours since 1992-1-1" ;

        double valtime(record) ;	// forecast time ("valid" time)
               valtime:long_name = "valid time" ;
               valtime:units = "hours since 1992-1-1" ;

        :record = "reftime, valtime" ;	// "dimension attribute" -- means
                                        // (reftime, valtime) uniquely
                                        // determine record

        char   datetime(record, time_len) ; // derived from reftime
               datetime:long_name = "reference date and time" ;
               // units YYYY-MM-DD hh:mm:ssZ  (ISO 8601)

        double valtime_offset(valtime_offset) ; // valtime - reftime
               valtime_offset:long_name = "hours from reference time" ;
               valtime_offset:units = "hours" ;

        char   forecasttime(record, time_len) ; // derived from valtime
               forecasttime:long_name = "forecast date and time" ;
               // units YYYY-MM-DD hh:mm:ssZ  (ISO 8601)

        float  level(level) ;
               level:long_name = "isobaric level" ;
               level:units = "hectopascals" ;


        // The following lat and lon coordinate variables are redundant,
        // since the navigation variables provide the necessary information.
        // The extra information is included here for human readability.

        float  lat(lat) ;
               lat:long_name = "latitude" ;
               lat:units = "degrees_north" ;

        float  lon(lon) ;
               lon:long_name = "longitude" ;
               lon:units = "degrees_east" ;

        long   model_id(nmodels) ;
               model_id:long_name = "generating process ID number" ;

        // navigation variables all use nav dimension

        char   nav_model(nav, nav_len) ;        // navigation parameterization
               nav_model:long_name = "navigation model name" ;

        int    grid_type_code(nav) ;
               grid_type_code:long_name = "GRIB-1 GDS data representation type" ;

        char   grid_type(nav, nav_len) ;
               grid_type:long_name = "GRIB-1 grid type" ;

        char   grid_name(nav, nav_len) ;
               grid_name:long_name = "grid name" ;

        int    grid_center(nav) ;
               grid_center:long_name = "GRIB-1 originating center ID" ;

        int    grid_number(nav, ngrids) ;
               grid_number:long_name = "GRIB-1 catalogued grid numbers" ;
               grid_number:_FillValue = -9999 ;

        char   i_dim(nav, nav_len) ;
               i_dim:long_name = "longitude dimension name" ;

        char   j_dim(nav, nav_len) ;
               j_dim:long_name = "latitude dimension name" ;

        int    Ni(nav) ;
               Ni:long_name = "number of points along a latitude circle" ;

        int    Nj(nav) ;
               Nj:long_name = "number of points along a longitude circle" ;

        float  La1(nav) ;
               La1:long_name = "latitude of first grid point" ;
               La1:units = "degrees_north" ;

        float  Lo1(nav) ;
               Lo1:long_name = "longitude of first grid point" ;
               Lo1:units = "degrees_east" ;

        float  La2(nav) ;
               La2:long_name = "latitude of last grid point" ;
               La2:units = "degrees_north" ;

        float  Lo2(nav) ;
               Lo2:long_name = "longitude of last grid point" ;
               Lo2:units = "degrees_east" ;

        float  Di(nav) ;
               Di:long_name = "longitudinal direction increment" ;
               Di:units = "degrees" ;

        float  Dj(nav) ;
               Dj:long_name = "latitudinal direction increment" ;
               Dj:units = "degrees" ;

        byte   ResCompFlag(nav) ;
               ResCompFlag:long_name = "resolution and component flags" ;

        // end of navigation variables

        float  P_msl(record,lat,lon) ;
               P_msl:long_name = "Pressure reduced to MSL at mean sea level" ;
               P_msl:standard_name = "air_pressure_at_sea_level" ;
               P_msl:units = "Pa" ;
               P_msl:GRIB_parameter_number = 2 ;
               P_msl:GRIB_level_flag = 102 ;
               P_msl:_FillValue = -9999.f ;
               P_msl:navigation = "nav" ;

        float  Z(record,level,lat,lon) ;
               Z:long_name = "Geopotential height at isobaric levels" ;
               Z:standard_name = "geopotential_height" ;
               Z:units = "gp m" ;
               Z:GRIB_parameter_number = 7 ;
               Z:GRIB_level_flag = 100 ;
               Z:_FillValue = -9999.f ;
               Z:navigation = "nav" ;

        float  u(record,level,lat,lon) ;
               u:long_name = "u-component of wind at isobaric levels" ;
               u:standard_name = "eastward_wind" ;
               u:units = "m/s" ;
               u:GRIB_parameter_number = 33 ;
               u:GRIB_level_flag = 100 ;
               u:_FillValue = -9999.f ;
               u:navigation = "nav" ;

        float  v(record,level,lat,lon) ;
               v:long_name = "v-component of wind at isobaric levels" ;
               v:standard_name = "northward_wind" ;
               v:units = "m/s" ;
               v:GRIB_parameter_number = 34 ;
               v:GRIB_level_flag = 100 ;
               v:_FillValue = -9999.f ;
               v:navigation = "nav" ;


// global attributes
               :history = "2003-04-04 14:44:21 - created by gribtocdl" ; 
               :title = "Medium Range Forecasts Extended" ;
               :Conventions = "NUWG" ;
               :GRIB_reference = "Office Note 388 GRIB" ;
               :GRIB_URL = "http://www.nco.ncep.noaa.gov/pmb/docs/on388/" ;
               :version = 1.0 ;

data:

 level = 1000.0, 500.0 ;
 model_id = 80, 94 ;
 valtime_offset = 84, 96, 108, 120, 132, 144, 156, 168, 180, 192, 204, 216, 228, 240 ;


 // Navigation
 nav_model = "GRIB1" ;
 grid_type_code = 0 ;
 grid_type = "Latitude/Longitude" ;
 grid_name = "Global 5.0 x 5.0 degree grid" ;
 grid_center = 7 ;
 grid_number = 25, 26 ;
 i_dim = "lon" ;
 j_dim = "lat" ;
 Ni = 72 ;
 Nj = 37 ;
 La1 = -90.000000 ;
 Lo1 = 0.000000 ;
 La2 = 90.000000 ;
 Lo2 = 355.000000 ;
 Di = 5.000000 ;
 Dj = 5.000000 ;
 ResCompFlag = 136 ;

 lon =  0.00,  5.00, 10.00, 15.00, 20.00, 25.00, 30.00, 35.00,
       40.00, 45.00, 50.00, 55.00, 60.00, 65.00, 70.00, 75.00,
       80.00, 85.00, 90.00, 95.00,100.00,105.00,110.00,115.00,
      120.00,125.00,130.00,135.00,140.00,145.00,150.00,155.00,
      160.00,165.00,170.00,175.00,180.00,185.00,190.00,195.00,
      200.00,205.00,210.00,215.00,220.00,225.00,230.00,235.00,
      240.00,245.00,250.00,255.00,260.00,265.00,270.00,275.00,
      280.00,285.00,290.00,295.00,300.00,305.00,310.00,315.00,
      320.00,325.00,330.00,335.00,340.00,345.00,350.00,355.00 ;

 lat =-90.00,-85.00,-80.00,-75.00,-70.00,-65.00,-60.00,-55.00,
      -50.00,-45.00,-40.00,-35.00,-30.00,-25.00,-20.00,-15.00,
      -10.00, -5.00,  0.00,  5.00, 10.00, 15.00, 20.00, 25.00,
       30.00, 35.00, 40.00, 45.00, 50.00, 55.00, 60.00, 65.00,
       70.00, 75.00, 80.00, 85.00, 90.00 ;

}
