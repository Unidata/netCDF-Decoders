netcdf eta{        // Early Terrain Analysis model 48km and 80km 

dimensions:
        record = UNLIMITED ;   // (reference time, forecast time)
        x = 93 ;
        y = 65 ;
        level = 19 ;           // isobaric levels
        alevel = 5 ;           // Absolute vorticity isobaric levels
        lpdg = 6 ;             // layer between levels at specif. pressure diffs from ground
        fhg = 2 ;              // fixed height above ground
        lfhg = 1 ;             // layer between 2 height levels above ground
        time_len = 21 ;        // string length for datetime strings
        valtime_offset = 11 ;  // number of offset times
        nmodels = 1 ;          // number of models
        ngrids = 1 ;           // number of grids
        nav = 1 ;              // for navigation
        nav_len = 100 ;        // max string length for navigation strings

variables:

        double reftime(record) ;	// reference time of the model
               reftime:long_name = "reference time" ;
               reftime:units = "hours since 1992-1-1" ;

        double valtime(record) ;	// forecast time ("valid" time)
               valtime:long_name = "valid time" ;
               valtime:units = "hours since 1992-1-1" ;

        :record = "reftime, valtime" ;	// "dimension attribute" -- means
                                        // (reftime, valtime) uniquely
                                        // determine record

        char   datetime(record, time_len) ; // derived from reftime
               datetime:long_name = "reference date and time" ;
               // units YYYY-MM-DD hh:mm:ssZ  (ISO 8601)

        double valtime_offset(valtime_offset) ; // valtime - reftime
               valtime_offset:long_name = "hours from reference time" ;
               valtime_offset:units = "hours" ;

        char   forecasttime(record, time_len) ; // derived from valtime
               forecasttime:long_name = "forecast date and time" ;
               // units YYYY-MM-DD hh:mm:ssZ  (ISO 8601)

        float  level(level) ;
               level:long_name = "isobaric level" ;
               level:units = "hectopascals" ;

        float  alevel(alevel) ;
               alevel:long_name = "isobaric level" ;
               alevel:units = "hectopascals" ;

        :lpdg = "lpdg_bot, lpdg_top" ; // ("lpdg_bot, lpdg_top") uniquely
                                       // determines lpdg

        float  lpdg_bot(lpdg) ;
               lpdg_bot:long_name = "bottom level of layer between levels at specif. pressure diffs from ground " ;
               lpdg_bot:units = "hPa" ;

        float  lpdg_top(lpdg) ;
               lpdg_top:long_name = "top level of layer between levels at specif. pressure diffs from ground " ;
               lpdg_top:units = "hPa" ;

        float  fhg(fhg) ;
               fhg:long_name = "fixed height above ground" ;
               fhg:units = "meters" ;

        :lfhg = "lfhg_bot, lfhg_top" ; // ("lfhg_bot, lfhg_top") uniquely
                                       // determines lfhg

        float  lfhg_bot(lfhg) ;
               lfhg_bot:long_name = "bottom level of layer between 2 height levels above ground " ;
               lfhg_bot:units = "hm" ;

        float  lfhg_top(lfhg) ;
               lfhg_top:long_name = "top level of layer between 2 height levels above ground " ;
               lfhg_top:units = "hm" ;


        long   model_id(nmodels) ;
               model_id:long_name = "generating process ID number" ;

        // navigation variables all use nav dimension

        char   nav_model(nav, nav_len) ;        // navigation parameterization
               nav_model:long_name = "navigation model name" ;

        int    grid_type_code(nav) ;
               grid_type_code:long_name = "GRIB-1 GDS data representation type" ;

        char   grid_type(nav, nav_len) ;
               grid_type:long_name = "GRIB-1 grid type" ;

        char   grid_name(nav, nav_len) ;
               grid_name:long_name = "grid name" ;

        int    grid_center(nav) ;
               grid_center:long_name = "GRIB-1 originating center ID" ;

        int    grid_number(nav, ngrids) ;
               grid_number:long_name = "GRIB-1 catalogued grid numbers" ;
               grid_number:_FillValue = -9999 ;

        char   x_dim(nav, nav_len) ;
               x_dim:long_name = "x dimension name" ;

        char   y_dim(nav, nav_len) ;
               y_dim:long_name = "y dimension name" ;

        long   Nx(nav) ;
               Nx:long_name = "number of points along x-axis" ;

        long   Ny(nav) ;
               Ny:long_name =  "number of points along y-axis" ;

        float  La1(nav) ;
               La1:long_name = "latitude of first grid point" ;
               La1:units = "degrees_north" ;

        float  Lo1(nav) ;
               Lo1:long_name = "longitude of first grid point" ;
               Lo1:units = "degrees_east" ;

        float  Lov(nav) ;
               Lov:long_name = "orientation of the grid" ;
               Lov:units = "degrees_east" ;

        float  Dx(nav) ;
               Dx:long_name = "x-direction grid length" ;
               Dx:units = "m" ;

        float  Dy(nav) ;
               Dy:long_name = "y-direction grid length" ;
               Dy:units = "m" ;

        byte   ProjFlag(nav) ;
               ProjFlag:long_name = "projection center flag" ;

        float  Latin1(nav) ;
               Latin1:long_name = "first intersecting latitude" ;
               Latin1:units = "degrees_north" ;

        float  Latin2(nav) ;
               Latin2:long_name = "second intersecting latitude" ;
               Latin2:units = "degrees_north" ;

        float  SpLat(nav) ;
               SpLat:long_name = "latitude of the southern pole" ;
               SpLat:units = "degrees_north" ;

        float  SpLon(nav) ;
               SpLon:long_name = "longitude of the southern pole" ;
               SpLon:units = "degrees_east" ;

        byte   ResCompFlag(nav) ;
               ResCompFlag:long_name = "resolution and component flags" ;

        // end of navigation variables

        float  omega(record,level,y,x) ;
               omega:long_name = "Pressure vertical velocity at isobaric levels" ;
               omega:standard_name = "omega" ;
               omega:units = "Pa/s" ;
               omega:GRIB_parameter_number = 39 ;
               omega:GRIB_level_flag = 100 ;
               omega:_FillValue = -9999.f ;
               omega:navigation = "nav" ;

        float  Z(record,level,y,x) ;
               Z:long_name = "Geopotential height at isobaric levels" ;
               Z:standard_name = "geopotential_height" ;
               Z:units = "gp m" ;
               Z:GRIB_parameter_number = 7 ;
               Z:GRIB_level_flag = 100 ;
               Z:_FillValue = -9999.f ;
               Z:navigation = "nav" ;

        float  Z_sfc(y,x) ;
               Z_sfc:long_name = "Geopotential height at surface of the earth" ;
               Z_sfc:standard_name = "geopotential_height" ;
               Z_sfc:units = "gp m" ;
               Z_sfc:GRIB_parameter_number = 7 ;
               Z_sfc:GRIB_level_flag = 1 ;
               Z_sfc:_FillValue = -9999.f ;
               Z_sfc:navigation = "nav" ;

        float  Z_frzlvl(record,y,x) ;
               Z_frzlvl:long_name = "Geopotential height at 0 degree isotherm level" ;
               Z_frzlvl:standard_name = "geopotential_height" ;
               Z_frzlvl:units = "gp m" ;
               Z_frzlvl:GRIB_parameter_number = 7 ;
               Z_frzlvl:GRIB_level_flag = 4 ;
               Z_frzlvl:_FillValue = -9999.f ;
               Z_frzlvl:navigation = "nav" ;

        float  v(record,level,y,x) ;
               v:long_name = "v-component of wind at isobaric levels" ;
               v:standard_name = "northward_wind" ;
               v:units = "m/s" ;
               v:GRIB_parameter_number = 34 ;
               v:GRIB_level_flag = 100 ;
               v:_FillValue = -9999.f ;
               v:navigation = "nav" ;

        float  v_fhg(record,fhg,y,x) ;
               v_fhg:long_name = "v-component of wind at fixed height above ground" ;
               v_fhg:standard_name = "northward_wind" ;
               v_fhg:units = "m/s" ;
               v_fhg:GRIB_parameter_number = 34 ;
               v_fhg:GRIB_level_flag = 105 ;
               v_fhg:_FillValue = -9999.f ;
               v_fhg:navigation = "nav" ;

        float  v_lpdg(record,lpdg,y,x) ;
               v_lpdg:long_name = "v-component of wind at layer between levels at specif. pressure diffs from ground" ;
               v_lpdg:standard_name = "northward_wind" ;
               v_lpdg:units = "m/s" ;
               v_lpdg:GRIB_parameter_number = 34 ;
               v_lpdg:GRIB_level_flag = 116 ;
               v_lpdg:_FillValue = -9999.f ;
               v_lpdg:navigation = "nav" ;

        float  v_trop(record,y,x) ;
               v_trop:long_name = "v-component of wind at tropopause" ;
               v_trop:standard_name = "northward_wind" ;
               v_trop:units = "m/s" ;
               v_trop:GRIB_parameter_number = 34 ;
               v_trop:GRIB_level_flag = 7 ;
               v_trop:_FillValue = -9999.f ;
               v_trop:navigation = "nav" ;

        float  v_maxwind(record,y,x) ;
               v_maxwind:long_name = "v-component of wind at maximium wind speed level" ;
               v_maxwind:standard_name = "northward_wind" ;
               v_maxwind:units = "m/s" ;
               v_maxwind:GRIB_parameter_number = 34 ;
               v_maxwind:GRIB_level_flag = 6 ;
               v_maxwind:_FillValue = -9999.f ;
               v_maxwind:navigation = "nav" ;

        float  T(record,level,y,x) ;
               T:long_name = "Temperature at isobaric levels" ;
               T:standard_name = "air_temperature" ;
               T:units = "degK" ;
               T:GRIB_parameter_number = 11 ;
               T:GRIB_level_flag = 100 ;
               T:_FillValue = -9999.f ;
               T:navigation = "nav" ;

        float  T_fhg(record,fhg,y,x) ;
               T_fhg:long_name = "Temperature at fixed height above ground" ;
               T_fhg:standard_name = "air_temperature" ;
               T_fhg:units = "degK" ;
               T_fhg:GRIB_parameter_number = 11 ;
               T_fhg:GRIB_level_flag = 105 ;
               T_fhg:_FillValue = -9999.f ;
               T_fhg:navigation = "nav" ;

        float  T_lpdg(record,lpdg,y,x) ;
               T_lpdg:long_name = "Temperature at layer between levels at specif. pressure diffs from ground" ;
               T_lpdg:standard_name = "air_temperature" ;
               T_lpdg:units = "degK" ;
               T_lpdg:GRIB_parameter_number = 11 ;
               T_lpdg:GRIB_level_flag = 116 ;
               T_lpdg:_FillValue = -9999.f ;
               T_lpdg:navigation = "nav" ;

        float  T_trop(record,y,x) ;
               T_trop:long_name = "Temperature at tropopause" ;
               T_trop:standard_name = "air_temperature" ;
               T_trop:units = "degK" ;
               T_trop:GRIB_parameter_number = 11 ;
               T_trop:GRIB_level_flag = 7 ;
               T_trop:_FillValue = -9999.f ;
               T_trop:navigation = "nav" ;

        float  T_cltp(record,y,x) ;
               T_cltp:long_name = "Temperature at cloud top level" ;
               T_cltp:standard_name = "air_temperature" ;
               T_cltp:GRIB_parameter_number = 11 ;
               T_cltp:GRIB_level_flag = 3 ;
               T_cltp:units = "degK" ;
               T_cltp:_FillValue = -9999.f ;
               T_cltp:navigation = "nav" ;

        float  u(record,level,y,x) ;
               u:long_name = "u-component of wind at isobaric levels" ;
               u:standard_name = "eastward_wind" ;
               u:units = "m/s" ;
               u:GRIB_parameter_number = 33 ;
               u:GRIB_level_flag = 100 ;
               u:_FillValue = -9999.f ;
               u:navigation = "nav" ;

        float  u_fhg(record,fhg,y,x) ;
               u_fhg:long_name = "u-component of wind at fixed height above ground" ;
               u_fhg:standard_name = "eastward_wind" ;
               u_fhg:units = "m/s" ;
               u_fhg:GRIB_parameter_number = 33 ;
               u_fhg:GRIB_level_flag = 105 ;
               u_fhg:_FillValue = -9999.f ;
               u_fhg:navigation = "nav" ;

        float  u_lpdg(record,lpdg,y,x) ;
               u_lpdg:long_name = "u-component of wind at layer between levels at specif. pressure diffs from ground" ;
               u_lpdg:standard_name = "eastward_wind" ;
               u_lpdg:units = "m/s" ;
               u_lpdg:GRIB_parameter_number = 33 ;
               u_lpdg:GRIB_level_flag = 116 ;
               u_lpdg:_FillValue = -9999.f ;
               u_lpdg:navigation = "nav" ;

        float  u_trop(record,y,x) ;
               u_trop:long_name = "u-component of wind at tropopause" ;
               u_trop:standard_name = "eastward_wind" ;
               u_trop:units = "m/s" ;
               u_trop:GRIB_parameter_number = 33 ;
               u_trop:GRIB_level_flag = 7 ;
               u_trop:_FillValue = -9999.f ;
               u_trop:navigation = "nav" ;

        float  u_maxwind(record,y,x) ;
               u_maxwind:long_name = "u-component of wind at maximium wind speed level" ;
               u_maxwind:standard_name = "eastward_wind" ;
               u_maxwind:units = "m/s" ;
               u_maxwind:GRIB_parameter_number = 33 ;
               u_maxwind:GRIB_level_flag = 6 ;
               u_maxwind:_FillValue = -9999.f ;
               u_maxwind:navigation = "nav" ;

        float  RH(record,level,y,x) ;
               RH:long_name = "Relative humidity at isobaric levels" ;
               RH:standard_name = "relative_humidity" ;
               RH:units = "percent" ;
               RH:GRIB_parameter_number = 52 ;
               RH:GRIB_level_flag = 100 ;
               RH:_FillValue = -9999.f ;
               RH:navigation = "nav" ;

        float  RH_fhg(record,fhg,y,x) ;
               RH_fhg:long_name = "Relative humidity at fixed height above ground" ;
               RH_fhg:standard_name = "relative_humidity" ;
               RH_fhg:units = "percent" ;
               RH_fhg:GRIB_parameter_number = 52 ;
               RH_fhg:GRIB_level_flag = 105 ;
               RH_fhg:_FillValue = -9999.f ;
               RH_fhg:navigation = "nav" ;

        float  RH_lpdg(record,lpdg,y,x) ;
               RH_lpdg:long_name = "Relative humidity at layer between levels at specif. pressure diffs from ground" ;
               RH_lpdg:standard_name = "relative_humidity" ;
               RH_lpdg:units = "percent" ;
               RH_lpdg:GRIB_parameter_number = 52 ;
               RH_lpdg:GRIB_level_flag = 116 ;
               RH_lpdg:_FillValue = -9999.f ;
               RH_lpdg:navigation = "nav" ;

        float  RH_frzlvl(record,y,x) ;
               RH_frzlvl:long_name = "Relative humidity at 0 degree isotherm level" ;
               RH_frzlvl:standard_name = "relative_humidity" ;
               RH_frzlvl:units = "percent" ;
               RH_frzlvl:GRIB_parameter_number = 52 ;
               RH_frzlvl:GRIB_level_flag = 4 ;
               RH_frzlvl:_FillValue = -9999.f ;
               RH_frzlvl:navigation = "nav" ;

        float  P_sfc(record,y,x) ;
               P_sfc:long_name = "Pressure at surface of the earth" ;
               P_sfc:standard_name = "air_pressure" ;
               P_sfc:units = "Pa" ;
               P_sfc:GRIB_parameter_number = 1 ;
               P_sfc:GRIB_level_flag = 1 ;
               P_sfc:_FillValue = -9999.f ;
               P_sfc:navigation = "nav" ;

        float  P_trop(record,y,x) ;
               P_trop:long_name = "Pressure at tropopause" ;
               P_trop:standard_name = "air_pressure" ;
               P_trop:units = "Pa" ;
               P_trop:GRIB_parameter_number = 1 ;
               P_trop:GRIB_level_flag = 7 ;
               P_trop:_FillValue = -9999.f ;
               P_trop:navigation = "nav" ;

        float  P_msl(record,y,x) ;
               P_msl:long_name = "Pressure reduced to MSL at mean sea level" ;
               P_msl:standard_name = "air_pressure_at_sea_level" ;
               P_msl:units = "Pa" ;
               P_msl:GRIB_parameter_number = 2 ;
               P_msl:GRIB_level_flag = 102 ;
               P_msl:_FillValue = -9999.f ;
               P_msl:navigation = "nav" ;

        float  P_maxwind(record,y,x) ;
               P_maxwind:long_name = "Pressure at maximium wind speed level" ;
               P_maxwind:standard_name = "air_pressure" ;
               P_maxwind:units = "Pa" ;
               P_maxwind:GRIB_parameter_number = 1 ;
               P_maxwind:GRIB_level_flag = 6 ;
               P_maxwind:_FillValue = -9999.f ;
               P_maxwind:navigation = "nav" ;

        float  P_clbs(record,y,x) ;
               P_clbs:long_name = "Pressure at cloud base level" ;
               P_clbs:standard_name = "air_pressure" ;
               P_clbs:GRIB_parameter_number = 1 ;
               P_clbs:GRIB_level_flag = 2 ;
               P_clbs:units = "Pa" ;
               P_clbs:_FillValue = -9999.f ;
               P_clbs:navigation = "nav" ;

        float  P_cltp(record,y,x) ;
               P_cltp:long_name = "Pressure at cloud top level" ;
               P_cltp:standard_name = "air_pressure" ;
               P_cltp:GRIB_parameter_number = 1 ;
               P_cltp:GRIB_level_flag = 3 ;
               P_cltp:units = "Pa" ;
               P_cltp:_FillValue = -9999.f ;
               P_cltp:navigation = "nav" ;

        float  PRECIP(record,y,x) ;
               PRECIP:long_name = "Total precipitation at surface of the earth" ;
               PRECIP:standard_name = "precipitation_amount" ;
               PRECIP:units = "kg/m2" ;
               PRECIP:GRIB_parameter_number = 61 ;
               PRECIP:GRIB_level_flag = 1 ;
               PRECIP:_FillValue = -9999.f ;
               PRECIP:navigation = "nav" ;

        float  precip_cn(record,y,x) ;
               precip_cn:long_name = "Convective precipitation at surface of the earth" ;
               precip_cn:standard_name = "convective_precipitation_amount" ;
               precip_cn:units = "kg/m2" ;
               precip_cn:GRIB_parameter_number = 63 ;
               precip_cn:GRIB_level_flag = 1 ;
               precip_cn:_FillValue = -9999.f ;
               precip_cn:navigation = "nav" ;

        float  Psl_et(record,y,x) ;
               Psl_et:long_name = "Mean sea level pressure (ETA model reduction) at mean sea level" ;
               Psl_et:standard_name = "-" ;
               Psl_et:units = "Pa" ;
               Psl_et:GRIB_parameter_number = 130 ;
               Psl_et:GRIB_level_flag = 102 ;
               Psl_et:_FillValue = -9999.f ;
               Psl_et:navigation = "nav" ;

        float  absvor(record,alevel,y,x) ;
               absvor:long_name = "Absolute vorticity at isobaric levels" ;
               absvor:standard_name = "atmosphere_absolute_vorticity" ;
               absvor:units = "1/s" ;
               absvor:GRIB_parameter_number = 41 ;
               absvor:GRIB_level_flag = 100 ;
               absvor:_FillValue = -9999.f ;
               absvor:navigation = "nav" ;

        float  pli_lpdg(record,lpdg,y,x) ;
               pli_lpdg:long_name = "Parcel lifted index (to 500 hPa) at layer between levels at specif. pressure diffs from ground" ;
               pli_lpdg:standard_name = "-" ;
               pli_lpdg:units = "K" ;
               pli_lpdg:GRIB_parameter_number = 24 ;
               pli_lpdg:GRIB_level_flag = 116 ;
               pli_lpdg:_FillValue = -9999.f ;
               pli_lpdg:navigation = "nav" ;

        float  LI4_lpdg(record,lpdg,y,x) ;
               LI4_lpdg:long_name = "Best (4 layer) lifted index at layer between levels at specif. pressure diffs from ground" ;
               LI4_lpdg:standard_name = "-" ;
               LI4_lpdg:units = "degK" ;
               LI4_lpdg:GRIB_parameter_number = 132 ;
               LI4_lpdg:GRIB_level_flag = 116 ;
               LI4_lpdg:_FillValue = -9999.f ;
               LI4_lpdg:navigation = "nav" ;

        float  pr_water_atm(record,y,x) ;
               pr_water_atm:long_name = "Precipitable water at entire atmosphere considered as a single layer" ;
               pr_water_atm:standard_name = "atmosphere_water_vapour_content" ;
               pr_water_atm:units = "kg/m2" ;
               pr_water_atm:GRIB_parameter_number = 54 ;
               pr_water_atm:GRIB_level_flag = 200 ;
               pr_water_atm:_FillValue = -9999.f ;
               pr_water_atm:navigation = "nav" ;

        float  cape_sfc(record,y,x) ;
               cape_sfc:long_name = "Convective available potential energy at surface of the earth" ;
               cape_sfc:standard_name = "-" ;
               cape_sfc:units = "J/kg" ;
               cape_sfc:GRIB_parameter_number = 157 ;
               cape_sfc:GRIB_level_flag = 1 ;
               cape_sfc:_FillValue = -9999.f ;
               cape_sfc:navigation = "nav" ;

        float  cape_lpdg(record,lpdg,y,x) ;
               cape_lpdg:long_name = "Convective available potential energy at layer between levels at specif. pressure diffs from ground" ;
               cape_lpdg:standard_name = "-" ;
               cape_lpdg:units = "J/kg" ;
               cape_lpdg:GRIB_parameter_number = 157 ;
               cape_lpdg:GRIB_level_flag = 116 ;
               cape_lpdg:_FillValue = -9999.f ;
               cape_lpdg:navigation = "nav" ;

        float  cin_lpdg(record,lpdg,y,x) ;
               cin_lpdg:long_name = "Convective inhibition at layer between levels at specif. pressure diffs from ground" ;
               cin_lpdg:standard_name = "-" ;
               cin_lpdg:units = "J/kg" ;
               cin_lpdg:GRIB_parameter_number = 156 ;
               cin_lpdg:GRIB_level_flag = 116 ;
               cin_lpdg:_FillValue = -9999.f ;
               cin_lpdg:navigation = "nav" ;

        float  cin_sfc(record,y,x) ;
               cin_sfc:long_name = "Convective inhibition at surface of the earth" ;
               cin_sfc:standard_name = "-" ;
               cin_sfc:units = "J/kg" ;
               cin_sfc:GRIB_parameter_number = 156 ;
               cin_sfc:GRIB_level_flag = 1 ;
               cin_sfc:_FillValue = -9999.f ;
               cin_sfc:navigation = "nav" ;

        float  helc_lfhg(record,lfhg,y,x) ;
               helc_lfhg:long_name = "Storm relative helicity at layer between 2 height levels above ground" ;
               helc_lfhg:standard_name = "-" ;
               helc_lfhg:units = "m2/s2" ;
               helc_lfhg:GRIB_parameter_number = 190 ;
               helc_lfhg:GRIB_level_flag = 106 ;
               helc_lfhg:_FillValue = -9999.f ;
               helc_lfhg:navigation = "nav" ;


// global attributes
               :history = "2003-03-28 11:00:39 - created by gribtocdl" ; 
               :title = " Early Terrain Analysis model 48km and 80km" ;
               :Conventions = "NUWG" ;
               :GRIB_reference = "Office Note 388 GRIB" ;
               :GRIB_URL = "http://www.nco.ncep.noaa.gov/pmb/docs/on388/" ;
               :version = 1.1 ;

data:

 level = 1000.0, 950.0, 900.0, 850.0, 800.0, 750.0, 700.0, 650.0, 600.0, 550.0, 
      500.0, 450.0, 400.0, 350.0, 300.0, 250.0, 200.0, 150.0, 100.0 ;
 alevel = 1000.0, 850.0, 700.0, 500.0, 250.0 ;
 lpdg_bot = 0.0, 0.0, 30.0, 60.0, 90.0, 120.0 ;
 lpdg_top = 30.0, 180.0, 60.0, 90.0, 120.0, 150.0 ;
 fhg = 2.0, 10.0 ;
 lfhg_bot = 0.0 ;
 lfhg_top = 30.0 ;
 model_id = 84 ;
 valtime_offset = 0, 6, 12, 18, 24, 30, 36, 42, 48, 54, 60 ;


 // Navigation
 nav_model = "GRIB1" ;
 grid_type_code = 3 ;
 grid_type = "Lambert conformal projection" ;
 grid_name = "grid 211: Regional CONUS" ;
 grid_center = 7 ;
 grid_number = 211 ;
 x_dim = "x" ;
 y_dim = "y" ;
 Nx = 93 ;
 Ny = 65 ;
 La1 = 12.190000 ;
 Lo1 = -133.459000 ;
 Lov = -95.000000 ;
 Dx = 81271.000000 ;
 Dy = 81271.000000 ;
 Latin1 = 25.000000 ;
 Latin2 = 25.000000 ;
 SpLat = 0.000000 ;
 SpLon = 0.000000 ;
 // Pole in proj. plane = North ;
 ProjFlag = 0 ;
 ResCompFlag = 8 ;

}
